library IEEE;
use IEEE.std_logic_1164.all;             -- Biblioteca para operações lógicas
use ieee.numeric_std.all;                -- Biblioteca para operações numéricas

-- Declaração da entidade memoriaROM com parâmetros genéricos para largura dos dados e endereços.
entity memoriaROM is
   generic (
          dataWidth: natural := 17;      -- Largura dos dados armazenados na memória
          addrWidth: natural := 9        -- Largura do endereço na memória
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);  -- Entrada de endereço
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)      -- Saída de dados
    );
end entity;

-- Arquitetura da memória ROM, nomeada como assincrona
architecture assincrona of memoriaROM is

  -- Tipo de dados para a memória, definido como um array de vetores lógicos.
  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);
  
  -- Definição das constantes para representar diferentes instruções.
  constant NOP   : std_logic_vector(3 downto 0) := "0000";
  constant LDA   : std_logic_vector(3 downto 0) := "0001";
  constant SOMA  : std_logic_vector(3 downto 0) := "0010";
  constant SUB   : std_logic_vector(3 downto 0) := "0011";
  constant LDI   : std_logic_vector(3 downto 0) := "0100";
  constant STA   : std_logic_vector(3 downto 0) := "0101";
  constant JMP   : std_logic_vector(3 downto 0) := "0110";
  constant JEQ   : std_logic_vector(3 downto 0) := "0111";
  constant CHECK : std_logic_vector(3 downto 0) := "1000";
  constant JSR   : std_logic_vector(3 downto 0) := "1001";
  constant RET   : std_logic_vector(3 downto 0) := "1010";
  constant ANDI  : std_logic_vector(3 downto 0) := "1011";
  constant JLT   : std_logic_vector(3 downto 0) := "1100";
  constant JNE   : std_logic_vector(3 downto 0) := "1101";
  
  -- Definição das constantes para os registros
  constant REG_0 : std_logic_vector(2 downto 0) := "000";
  constant REG_1 : std_logic_vector(2 downto 0) := "001";
  constant REG_2 : std_logic_vector(2 downto 0) := "010";
  constant REG_3 : std_logic_vector(2 downto 0) := "011";
  constant REG_4 : std_logic_vector(2 downto 0) := "100";
  constant REG_5 : std_logic_vector(2 downto 0) := "101";
  constant REG_6 : std_logic_vector(2 downto 0) := "110";
  constant REG_7 : std_logic_vector(2 downto 0) := "111";

  -- Função para inicializar a memória com instruções pré-definidas.
  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin

    -- Configurações de dados na memória
  
tmp(0) := LDI & REG_0 & "0000000000"; --  Inicializa R0 com 0
tmp(1) := LDI & REG_1 & "0000000001"; --  Inicializa R1 com 1
tmp(2) := LDI & REG_2 & "0000001010"; --  Inicializa R2 com 10
tmp(3) := LDI & REG_3 & "0000000110"; --  Inicializa R3 com 60
tmp(4) := LDI & REG_4 & "0000000010"; --  Inicializa R4 com 2
tmp(5) := LDI & REG_5 & "0000000100"; --  Inicializa R5 com 4
tmp(6) := LDI & REG_6 & "0010000000"; --  Inicializa R6 com 128
tmp(7) := LDI & REG_7 & "0000000011"; --  Inicializa R7 com 3
tmp(8) := STA & REG_0 & "0100100000"; --  0 -> HEX0
tmp(9) := STA & REG_0 & "0100100001"; --  0 -> HEX1
tmp(10) := STA & REG_0 & "0100100010"; --  0 -> HEX2
tmp(11) := STA & REG_0 & "0100100011"; --  0 -> HEX3
tmp(12) := STA & REG_0 & "0100100100"; --  0 -> HEX4
tmp(13) := STA & REG_0 & "0100100101"; --  0 -> HEX5
tmp(14) := STA & REG_0 & "0100000000"; --  0 -> LEDR0 ~ LEDR7
tmp(15) := STA & REG_0 & "0100000001"; --  0 -> LEDR8
tmp(16) := STA & REG_0 & "0100000010"; --  0 -> LEDR9
tmp(17) := STA & REG_0 & "0000000000"; --  0 -> Valor das unidades dos segundos
tmp(18) := STA & REG_0 & "0000000001"; --  0 -> Valor das dezenas dos segundos
tmp(19) := STA & REG_0 & "0000000010"; --  0 -> Valor das unidades dos minutos
tmp(20) := STA & REG_0 & "0000000011"; --  0 -> Valor das dezenas dos minutos
tmp(21) := STA & REG_0 & "0000000100"; --  0 -> Valor das unidades das horas
tmp(22) := STA & REG_0 & "0000000101"; --  0 -> Valor das dezenas das horas
tmp(23) := STA & REG_0 & "0000000110"; -- STA
tmp(24) := STA & REG_1 & "0000000111"; -- STA
tmp(25) := STA & REG_2 & "0000001000"; -- STA
tmp(26) := STA & REG_3 & "0000001001"; -- STA
tmp(27) := STA & REG_4 & "0000001010"; -- STA
tmp(28) := STA & REG_5 & "0000001011"; -- STA
tmp(29) := STA & REG_6 & "0000001100"; -- STA
tmp(30) := STA & REG_7 & "0000001101"; -- STA
tmp(31) := STA & REG_0 & "0000001110"; -- STA
tmp(32) := STA & REG_0 & "0000001111"; --  0 -> Novo valor das unidades dos segundos do alarme
tmp(33) := STA & REG_0 & "0000010000"; --  0 -> Novo valor das dezenas dos segundos do alarme
tmp(34) := STA & REG_0 & "0000010001"; --  0 -> Novo valor das unidades dos minutos do alarme
tmp(35) := STA & REG_0 & "0000010010"; --  0 -> Novo valor das dezenas dos minutos do alarme
tmp(36) := STA & REG_0 & "0000010011"; --  0 -> Novo valor das unidades das horas do alarme
tmp(37) := STA & REG_0 & "0000010100"; --  0 -> Novo valor das dezenas das horas do alarme
tmp(38) := STA & REG_0 & "0000010101"; --  0 -> Novo valor das unidades dos segundos
tmp(39) := STA & REG_0 & "0000010110"; --  0 -> Novo valor das dezenas dos segundos
tmp(40) := STA & REG_0 & "0000010111"; --  0 -> Novo valor das unidades dos minutos
tmp(41) := STA & REG_0 & "0000011000"; --  0 -> Novo valor das dezenas dos minutos
tmp(42) := STA & REG_0 & "0000011001"; --  0 -> Novo valor das unidades das horas
tmp(43) := STA & REG_0 & "0000011010"; --  0 -> Novo valor das dezenas das horas
tmp(44) := STA & REG_0 & "0000011011"; --  0 -> Flag timer
tmp(45) := STA & REG_0 & "0000011100"; --  0 -> Flag de ajuste das unidades dos segundos do timer
tmp(46) := STA & REG_0 & "0000011101"; --  0 -> Flag de ajuste das dezenas dos segundos do timer
tmp(47) := STA & REG_0 & "0000011110"; --  0 -> Flag de ajuste das unidades dos minutos do timer
tmp(48) := STA & REG_0 & "0000011111"; --  0 -> Flag de ajuste das dezenas dos minutos do timer
tmp(49) := STA & REG_0 & "0000100000"; --  0 -> Flag de ajuste das unidades das horas do timer
tmp(50) := STA & REG_0 & "0000100001"; --  0 -> Flag de ajuste das dezenas (>= 2) das horas do timer
tmp(51) := STA & REG_0 & "0000100010"; --  0 -> Flag de ajuste das dezenas (< 2) das horas do timer
tmp(52) := LDI & REG_3 & "0011111111"; -- LDI
tmp(53) := STA & REG_3 & "0000100011"; -- STA
tmp(54) := STA & REG_0 & "0000100100"; --  0 -> Flag de timer finalizado
tmp(55) := STA & REG_0 & "0000100101"; --  0 -> Flag de ajuste das unidades dos segundos do alarme
tmp(56) := STA & REG_0 & "0000100110"; --  0 -> Flag de ajuste das dezenas dos segundos do alarme
tmp(57) := STA & REG_0 & "0000100111"; --  0 -> Flag de ajuste das unidades dos minutos do alarme
tmp(58) := STA & REG_0 & "0000101000"; --  0 -> Flag de ajuste das dezenas dos minutos do alarme
tmp(59) := STA & REG_0 & "0000101001"; --  0 -> Flag de ajuste das unidades das horas do alarme
tmp(60) := STA & REG_0 & "0000101010"; --  0 -> Flag de ajuste das dezenas (>= 2) das horas do alarme
tmp(61) := STA & REG_0 & "0000101011"; --  0 -> Flag de ajuste das dezenas (< 2) das horas do alarme
tmp(62) := STA & REG_0 & "0000101100"; --  0 -> Flag de chegou no horário do alarme
tmp(63) := LDI & REG_3 & "0000001111"; -- LDI
tmp(64) := STA & REG_3 & "0000101101"; -- STA
tmp(65) := LDI & REG_3 & "0001000000"; -- LDI
tmp(66) := STA & REG_3 & "0000101110"; -- STA
tmp(67) := STA & REG_0 & "0111111111"; -- STA
tmp(68) := STA & REG_0 & "0111111110"; -- STA
tmp(69) := STA & REG_0 & "0111111101"; -- STA
tmp(70) := STA & REG_0 & "0111111100"; -- STA
tmp(71) := STA & REG_0 & "0111111011"; -- STA
tmp(72) := JSR & REG_0 & "0010110000"; -- JSR
tmp(73) := JSR & REG_0 & "0110110000"; -- JSR
tmp(74) := JSR & REG_0 & "0101101100"; -- JSR
tmp(75) := JSR & REG_0 & "0110001000"; -- JSR
tmp(76) := JSR & REG_0 & "0110011100"; -- JSR
tmp(77) := JSR & REG_0 & "1000101001"; -- JSR
tmp(78) := JSR & REG_0 & "0010010010"; -- JSR
tmp(79) := LDA & REG_6 & "0101100100"; --  Carrega o valor do Time Counter para R6
tmp(80) := ANDI & REG_6 & "0000000111"; -- ANDI
tmp(81) := CHECK & REG_6 & "0000000111"; --  Verifica se o Time Counter é igual a 0
tmp(82) := JNE & REG_0 & "0001001000"; -- JNE
tmp(83) := JSR & REG_0 & "0001010111"; -- JSR
tmp(84) := JSR & REG_0 & "0100100110"; -- JSR
tmp(85) := STA & REG_0 & "0111111011"; --  Limpa Leitura do Time Counter
tmp(86) := JMP & REG_0 & "0001001000"; -- JMP
tmp(87) := LDA & REG_7 & "0000000000"; --  Carrega o valor das unidades dos segundos para R7
tmp(88) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das unidades dos segundos
tmp(89) := STA & REG_7 & "0000000000"; --  Salva o valor das unidades dos segundos
tmp(90) := LDA & REG_7 & "0000000000"; --  Carrega o valor das unidades dos segundos para R7
tmp(91) := CHECK & REG_7 & "0000001000"; --  Verifica se o valor das unidades dos segundos é igual a 10
tmp(92) := JNE & REG_0 & "1001100001"; -- JNE
tmp(93) := STA & REG_0 & "0000000000"; --  0 -> Valor das unidades dos segundos
tmp(94) := LDA & REG_7 & "0000000001"; --  Carrega o valor das dezenas dos segundos para R7
tmp(95) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das dezenas dos segundos
tmp(96) := STA & REG_7 & "0000000001"; --  Salva o valor das dezenas dos segundos
tmp(97) := LDA & REG_7 & "0000000001"; --  Carrega o valor das dezenas dos segundos para R7
tmp(98) := CHECK & REG_7 & "0000001001"; --  Verifica se o valor das dezenas dos segundos é igual a 6
tmp(99) := JNE & REG_0 & "1001100001"; -- JNE
tmp(100) := STA & REG_0 & "0000000001"; --  0 -> Valor das dezenas dos segundos
tmp(101) := LDA & REG_7 & "0000000010"; --  Carrega o valor das unidades dos minutos para R7
tmp(102) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das unidades dos minutos
tmp(103) := STA & REG_7 & "0000000010"; --  Salva o valor das unidades dos minutos
tmp(104) := LDA & REG_7 & "0000000010"; --  Carrega o valor das unidades dos minutos para R7
tmp(105) := CHECK & REG_7 & "0000001000"; --  Verifica se o valor das unidades dos minutos é igual a 10
tmp(106) := JNE & REG_0 & "1001100001"; -- JNE
tmp(107) := STA & REG_0 & "0000000010"; --  0 -> Valor das unidades dos minutos
tmp(108) := LDA & REG_7 & "0000000011"; --  Carrega o valor das dezenas dos minutos para R7
tmp(109) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das dezenas dos minutos
tmp(110) := STA & REG_7 & "0000000011"; --  Salva o valor das dezenas dos minutos
tmp(111) := LDA & REG_7 & "0000000011"; --  Carrega o valor das dezenas dos minutos para R7
tmp(112) := CHECK & REG_7 & "0000001001"; --  Verifica se o valor das dezenas dos minutos é igual a 6
tmp(113) := JNE & REG_0 & "1001100001"; -- JNE
tmp(114) := STA & REG_0 & "0000000011"; --  0 -> Valor das dezenas dos minutos
tmp(115) := JSR & REG_0 & "0001110101"; -- JSR
tmp(116) := JMP & REG_0 & "1001100001"; -- JMP
tmp(117) := LDA & REG_7 & "0000000101"; --  Carrega o valor das dezenas das horas para R7
tmp(118) := CHECK & REG_7 & "0000001010"; --  Verifica se o valor das dezenas dos minutos é igual a 2
tmp(119) := JEQ & REG_0 & "0010000011"; -- JEQ
tmp(120) := LDA & REG_7 & "0000000100"; --  Carrega o valor das unidades das horas para R7
tmp(121) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das unidades das horas
tmp(122) := STA & REG_7 & "0000000100"; --  Salva o valor das unidades das horas
tmp(123) := LDA & REG_7 & "0000000100"; --  Carrega o valor das unidades das horas para R7
tmp(124) := CHECK & REG_7 & "0000001000"; --  Verifica se o valor das unidades das horas é igual a 10
tmp(125) := JNE & REG_0 & "1001100001"; -- JNE
tmp(126) := STA & REG_0 & "0000000100"; --  0 -> Valor das unidades das horas
tmp(127) := LDA & REG_7 & "0000000101"; --  Carrega o valor das dezenas das horas para R7
tmp(128) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das dezenas das horas
tmp(129) := STA & REG_7 & "0000000101"; --  Salva o valor das dezenas das horas
tmp(130) := RET & REG_0 & "0000000000"; -- RET
tmp(131) := LDA & REG_7 & "0000000100"; --  Carrega o valor das unidades das horas para R7
tmp(132) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das unidades das horas
tmp(133) := STA & REG_7 & "0000000100"; --  Salva o valor das unidades das horas
tmp(134) := LDA & REG_7 & "0000000100"; --  Carrega o valor das unidades das horas para R7
tmp(135) := CHECK & REG_7 & "0000001011"; --  Verifica se o valor das unidades das horas é igual a 4
tmp(136) := JNE & REG_0 & "1001100001"; -- JNE
tmp(137) := STA & REG_0 & "0000000100"; --  0 -> Valor das unidades das horas
tmp(138) := LDA & REG_7 & "0000000101"; --  Carrega o valor das dezenas das horas para R7
tmp(139) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das dezenas das horas
tmp(140) := STA & REG_7 & "0000000101"; --  Salva o valor das dezenas das horas
tmp(141) := LDA & REG_7 & "0000000101"; --  Carrega o valor das dezenas das horas para R7
tmp(142) := CHECK & REG_7 & "0000001101"; --  Verifica se o valor das dezenas das horas é igual a 3
tmp(143) := JNE & REG_0 & "1001100001"; -- JNE
tmp(144) := STA & REG_0 & "0000000101"; --  0 -> Valor das dezenas das horas
tmp(145) := RET & REG_0 & "0000000000"; -- RET
tmp(146) := LDA & REG_7 & "0101000000"; --  Carrega o valor dos SW0 até SW7 para R7
tmp(147) := ANDI & REG_7 & "0000101110"; --  Aplica máscara AND para isolar o bit 6
tmp(148) := CHECK & REG_7 & "0000101110"; --  Verifica se o bit 6 está setado
tmp(149) := JEQ & REG_0 & "0010100011"; -- JEQ
tmp(150) := LDA & REG_7 & "0000000101"; --  Carrega o valor das dezenas das horas para R7
tmp(151) := STA & REG_7 & "0100100101"; --  Salva o valor das dezenas das horas em HEX5
tmp(152) := LDA & REG_7 & "0000000100"; --  Carrega o valor das unidades das horas para R7
tmp(153) := STA & REG_7 & "0100100100"; --  Salva o valor das unidades das horas em HEX4
tmp(154) := LDA & REG_7 & "0000000011"; --  Carrega o valor das dezenas dos minutos para R7
tmp(155) := STA & REG_7 & "0100100011"; --  Salva o valor das dezenas dos minutos em HEX3
tmp(156) := LDA & REG_7 & "0000000010"; --  Carrega o valor das unidades dos minutos para R7
tmp(157) := STA & REG_7 & "0100100010"; --  Salva o valor das unidades dos minutos em HEX2
tmp(158) := LDA & REG_7 & "0000000001"; --  Carrega o valor das dezenas dos segundos para R7
tmp(159) := STA & REG_7 & "0100100001"; --  Salva o valor das dezenas dos segundos em HEX1
tmp(160) := LDA & REG_7 & "0000000000"; --  Carrega o valor das unidades dos segundos para R7
tmp(161) := STA & REG_7 & "0100100000"; --  Salva o valor das unidades dos segundos em HEX0
tmp(162) := RET & REG_0 & "0000000000"; -- RET
tmp(163) := LDA & REG_7 & "0000011010"; --  Carrega o valor das dezenas das horas do timer para R7
tmp(164) := STA & REG_7 & "0100100101"; --  Salva o valor das dezenas das horas do timer em HEX5
tmp(165) := LDA & REG_7 & "0000011001"; --  Carrega o valor das unidades das horas do timer para R7
tmp(166) := STA & REG_7 & "0100100100"; --  Salva o valor das unidades das horas do timer em HEX4
tmp(167) := LDA & REG_7 & "0000011000"; --  Carrega o valor das dezenas dos minutos do timer para R7
tmp(168) := STA & REG_7 & "0100100011"; --  Salva o valor das dezenas dos minutos do timer em HEX3
tmp(169) := LDA & REG_7 & "0000010111"; --  Carrega o valor das unidades dos minutos do timer para R7
tmp(170) := STA & REG_7 & "0100100010"; --  Salva o valor das unidades dos minutos do timer em HEX2
tmp(171) := LDA & REG_7 & "0000010110"; --  Carrega o valor das dezenas dos segundos do timer para R7
tmp(172) := STA & REG_7 & "0100100001"; --  Salva o valor das dezenas dos segundos do timer em HEX1
tmp(173) := LDA & REG_7 & "0000010101"; --  Carrega o valor das unidades dos segundos do timer para R7
tmp(174) := STA & REG_7 & "0100100000"; --  Salva o valor das unidades dos segundos do timer em HEX0
tmp(175) := RET & REG_0 & "0000000000"; -- RET
tmp(176) := LDA & REG_7 & "0101000000"; --  Carrega o R7 com a leitura das chaves SW0 até SW7
tmp(177) := ANDI & REG_7 & "0000001100"; --  Aplica máscara AND para isolar o bit 7
tmp(178) := CHECK & REG_7 & "0000001100"; --  Verifica se a chave SW7 está pressionada
tmp(179) := JEQ & REG_0 & "1001100001"; -- JEQ
tmp(180) := LDA & REG_7 & "0101100000"; --  Carrega o valor do botão KEY0
tmp(181) := ANDI & REG_7 & "0000000111"; --  Aplica máscara AND para isolar o bit 0
tmp(182) := CHECK & REG_7 & "0000000111"; --  Se KEY0 estiver pressionada, passa a setar o limite de incremento
tmp(183) := STA & REG_0 & "0111111111"; -- STA
tmp(184) := JNE & REG_0 & "1001100001"; -- JNE
tmp(185) := LDA & REG_7 & "0000011011"; --  Carrega o valor da flag de timer para R7
tmp(186) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de timer está setada
tmp(187) := JEQ & REG_0 & "1001100001"; -- JEQ
tmp(188) := STA & REG_1 & "0100000001"; --  Acende o LEDR8 para indicar que é o timer que está sendo setado, e não o alarme
tmp(189) := JSR & REG_0 & "1001011011"; -- JSR
tmp(190) := LDA & REG_7 & "0000100010"; --  Carrega o valor da flag de ajuste das dezenas (< 2) das horas para R7
tmp(191) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das dezenas das horas está setada
tmp(192) := JEQ & REG_0 & "0011010000"; -- JEQ
tmp(193) := LDA & REG_7 & "0000100001"; --  Carrega o valor da flag de ajuste das dezenas (>= 2) das horas para R7
tmp(194) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das dezenas das horas está setada
tmp(195) := JEQ & REG_0 & "0011011110"; -- JEQ
tmp(196) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(197) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(198) := STA & REG_7 & "0000011010"; --  Salva o valor de SW0 até SW7 em @26
tmp(199) := LDA & REG_7 & "0000011010"; --  Carrega o valor de SW0 até SW7 para R7
tmp(200) := CHECK & REG_7 & "0000001010"; --  Compara o valor de SW0 até SW7 com 2
tmp(201) := JLT & REG_0 & "0011001100"; -- JLT
tmp(202) := JEQ & REG_0 & "0011011010"; -- JEQ
tmp(203) := JMP & REG_0 & "1001100001"; -- JMP
tmp(204) := LDI & REG_3 & "0000100000"; --  Seta o valor 32 para R3
tmp(205) := STA & REG_3 & "0100000000"; --  Acende o LEDR5 para indicar que o valor das dezenas das horas do timer foi setado
tmp(206) := STA & REG_1 & "0000100010"; --  Ativa a flag de ajuste das dezenas das horas
tmp(207) := RET & REG_0 & "0000000000"; -- RET
tmp(208) := LDA & REG_7 & "0000100000"; --  Carrega o valor da flag de ajuste das unidades das horas para R7
tmp(209) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das unidades das horas está setada
tmp(210) := JEQ & REG_0 & "0011101100"; -- JEQ
tmp(211) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(212) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(213) := STA & REG_7 & "0000011001"; --  Salva o valor de SW0 até SW7 em @25
tmp(214) := LDA & REG_7 & "0000011001"; --  Carrega o valor de SW0 até SW7 para R7
tmp(215) := CHECK & REG_7 & "0000001000"; --  Compara o valor de SW0 até SW7 com 10
tmp(216) := JLT & REG_0 & "0011101000"; -- JLT
tmp(217) := JMP & REG_0 & "1001100001"; -- JMP
tmp(218) := LDI & REG_3 & "0000100000"; --  Seta o valor 32 para R3
tmp(219) := STA & REG_3 & "0100000000"; --  Acende o LEDR5 para indicar que o valor das dezenas das horas do timer foi setado
tmp(220) := STA & REG_1 & "0000100001"; --  Ativa a flag de ajuste das dezenas das horas
tmp(221) := RET & REG_0 & "0000000000"; -- RET
tmp(222) := LDA & REG_7 & "0000100000"; --  Carrega o valor da flag de ajuste das unidades das horas para R7
tmp(223) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das unidades das horas está setada
tmp(224) := JEQ & REG_0 & "0011101100"; -- JEQ
tmp(225) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(226) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(227) := STA & REG_7 & "0000011001"; --  Salva o valor de SW0 até SW7 em @25
tmp(228) := LDA & REG_7 & "0000011001"; --  Carrega o valor de SW0 até SW7 para R7
tmp(229) := CHECK & REG_7 & "0000001011"; --  Compara o valor de SW0 até SW7 com 4
tmp(230) := JLT & REG_0 & "0011101000"; -- JLT
tmp(231) := JMP & REG_0 & "1001100001"; -- JMP
tmp(232) := LDI & REG_3 & "0000110000"; --  Seta o valor 48 para R3
tmp(233) := STA & REG_3 & "0100000000"; --  Acende o LEDR5 e LEDR4 para indicar que os valores das dezenas e unidade de horas do timer foram setados
tmp(234) := STA & REG_1 & "0000100000"; --  Ativa a flag de ajuste das unidades das horas
tmp(235) := RET & REG_0 & "0000000000"; -- RET
tmp(236) := LDA & REG_7 & "0000011111"; --  Carrega o valor da flag de ajuste das dezenas dos minutos para R7
tmp(237) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das dezenas dos minutos está setada
tmp(238) := JEQ & REG_0 & "0011111010"; -- JEQ
tmp(239) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(240) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(241) := STA & REG_7 & "0000011000"; --  Salva o valor de SW0 até SW7 em @24
tmp(242) := LDA & REG_7 & "0000011000"; --  Carrega o valor de SW0 até SW7 para R7
tmp(243) := CHECK & REG_7 & "0000001001"; --  Compara o valor de SW0 até SW7 com 6
tmp(244) := JLT & REG_0 & "0011110110"; -- JLT
tmp(245) := JMP & REG_0 & "1001100001"; -- JMP
tmp(246) := LDI & REG_3 & "0000111000"; --  Seta o valor 56 para R3
tmp(247) := STA & REG_3 & "0100000000"; --  Acende o LEDR5, LEDR4 e LEDR3 para indicar que os valores das dezenas, unidade de horas e dezenas de minutos do timer foram setados
tmp(248) := STA & REG_1 & "0000011111"; --  Ativa a flag de ajuste das dezenas dos minutos
tmp(249) := RET & REG_0 & "0000000000"; -- RET
tmp(250) := LDA & REG_7 & "0000011110"; --  Carrega o valor da flag de ajuste das unidades dos minutos para R7
tmp(251) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das unidades dos minutos está setada
tmp(252) := JEQ & REG_0 & "0100001000"; -- JEQ
tmp(253) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(254) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(255) := STA & REG_7 & "0000010111"; --  Salva o valor de SW0 até SW7 em @23
tmp(256) := LDA & REG_7 & "0000010111"; --  Carrega o valor de SW0 até SW7 para R7
tmp(257) := CHECK & REG_7 & "0000001000"; --  Compara o valor de SW0 até SW7 com 10
tmp(258) := JLT & REG_0 & "0100000100"; -- JLT
tmp(259) := JMP & REG_0 & "1001100001"; -- JMP
tmp(260) := LDI & REG_3 & "0000111100"; --  Seta o valor 60 para R3
tmp(261) := STA & REG_3 & "0100000000"; --  Acende os LEDR5, LEDR4, LEDR3 e LEDR2 para indicar que os valores das dezenas, unidade de horas e dezenas de minutos do timer foram setados
tmp(262) := STA & REG_1 & "0000011110"; --  Ativa a flag de ajuste das unidades dos minutos
tmp(263) := RET & REG_0 & "0000000000"; -- RET
tmp(264) := LDA & REG_7 & "0000011101"; --  Carrega o valor da flag de ajuste das dezenas dos segundos para R7
tmp(265) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das dezenas dos segundos está setada
tmp(266) := JEQ & REG_0 & "0100010110"; -- JEQ
tmp(267) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(268) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(269) := STA & REG_7 & "0000010110"; --  Salva o valor de SW0 até SW7 em @22
tmp(270) := LDA & REG_7 & "0000010110"; --  Carrega o valor de SW0 até SW7 para R7
tmp(271) := CHECK & REG_7 & "0000001001"; --  Compara o valor de SW0 até SW7 com 6
tmp(272) := JLT & REG_0 & "0100010010"; -- JLT
tmp(273) := JMP & REG_0 & "1001100001"; -- JMP
tmp(274) := LDI & REG_3 & "0000111110"; --  Seta o valor 62 para R3
tmp(275) := STA & REG_3 & "0100000000"; --  Acende o LEDR5, LEDR4, LEDR3, LEDR2 e LEDR1 para indicar que os valores das dezenas, unidade de horas, dezenas e unidade de minutos e dezenas dos segundos do timer foram setados
tmp(276) := STA & REG_1 & "0000011101"; --  Ativa a flag de ajuste das dezenas dos segundos
tmp(277) := RET & REG_0 & "0000000000"; -- RET
tmp(278) := LDA & REG_7 & "0000011100"; --  Carrega o valor da flag de ajuste das unidades dos segundos para R7
tmp(279) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das unidades dos segundos está setada
tmp(280) := JEQ & REG_0 & "0100100000"; -- JEQ
tmp(281) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(282) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(283) := STA & REG_7 & "0000010101"; --  Salva o valor de SW0 até SW7 em @21
tmp(284) := LDA & REG_7 & "0000010101"; --  Carrega o valor de SW0 até SW7 para R7
tmp(285) := CHECK & REG_7 & "0000001000"; --  Compara o valor de SW0 até SW7 com 10
tmp(286) := JLT & REG_0 & "0100100000"; -- JLT
tmp(287) := JMP & REG_0 & "1001100001"; -- JMP
tmp(288) := LDI & REG_3 & "0000111111"; --  Seta o valor 63 para R3
tmp(289) := STA & REG_3 & "0100000000"; --  Acende o LEDR5, LEDR4, LEDR3, LEDR2, LEDR1 e LEDR0 para indicar que os valores das dezenas, unidade de horas, dezenas e unidade de minutos e dezenas e unidade dos segundos do timer foram setados
tmp(290) := STA & REG_1 & "0000011100"; --  Ativa a flag de ajuste das unidades dos segundos
tmp(291) := STA & REG_1 & "0000011011"; --  Ativa a flag de timer setado
tmp(292) := STA & REG_0 & "0000100100"; --  0 -> Flag de timer finalizado
tmp(293) := RET & REG_0 & "0000000000"; -- RET
tmp(294) := LDA & REG_7 & "0000011011"; --  Carrega o valor da flag de timer para R7
tmp(295) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de timer está setada
tmp(296) := JNE & REG_0 & "1001100001"; -- JNE
tmp(297) := LDA & REG_7 & "0000100100"; --  Carrega o valor da flag de timer finalizado para R7
tmp(298) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de timer finalizado está setada
tmp(299) := JEQ & REG_0 & "1001100001"; -- JEQ
tmp(300) := LDA & REG_7 & "0000010101"; --  Carrega o valor das unidades dos segundos do timer para R7
tmp(301) := SUB & REG_7 & "0000000111"; --  Decrementa o valor das unidades dos segundos do timer
tmp(302) := STA & REG_7 & "0000010101"; --  Salva o valor das unidades dos segundos do timer
tmp(303) := LDA & REG_7 & "0000100011"; --  Carrega o valor -1 para R7
tmp(304) := CHECK & REG_7 & "0000010101"; --  Verifica se o valor das unidades dos segundos do timer é igual a -1
tmp(305) := JNE & REG_0 & "1001100001"; -- JNE
tmp(306) := LDI & REG_3 & "0000001001"; --  Seta o valor 9 para R3
tmp(307) := STA & REG_3 & "0000010101"; --  Salva o valor 9 nas unidades dos segundos do timer
tmp(308) := LDA & REG_7 & "0000010110"; --  Carrega o valor das dezenas dos segundos do timer para R7
tmp(309) := SUB & REG_7 & "0000000111"; --  Decrementa o valor das dezenas dos segundos do timer
tmp(310) := STA & REG_7 & "0000010110"; --  Salva o valor das dezenas dos segundos do timer
tmp(311) := LDA & REG_7 & "0000100011"; --  Carrega o valor -1 para R7
tmp(312) := CHECK & REG_7 & "0000010110"; --  Verifica se o valor das dezenas dos segundos do timer é igual a -1
tmp(313) := JNE & REG_0 & "1001100001"; -- JNE
tmp(314) := LDI & REG_3 & "0000000101"; --  Seta o valor 5 para R3
tmp(315) := STA & REG_3 & "0000010110"; --  Salva o valor 5 nas dezenas dos segundos do timer
tmp(316) := LDA & REG_7 & "0000010111"; --  Carrega o valor das unidades dos minutos do timer para R7
tmp(317) := SUB & REG_7 & "0000000111"; --  Decrementa o valor das unidades dos minutos do timer
tmp(318) := STA & REG_7 & "0000010111"; --  Salva o valor das unidades dos minutos do timer
tmp(319) := LDA & REG_7 & "0000100011"; --  Carrega o valor -1 para R7
tmp(320) := CHECK & REG_7 & "0000010111"; --  Verifica se o valor das unidades dos minutos do timer é igual a -1
tmp(321) := JNE & REG_0 & "1001100001"; -- JNE
tmp(322) := LDI & REG_3 & "0000001001"; --  Seta o valor 9 para R3
tmp(323) := STA & REG_3 & "0000010111"; --  Salva o valor 9 nas unidades dos minutos do timer
tmp(324) := LDA & REG_7 & "0000011000"; --  Carrega o valor das dezenas dos minutos do timer para R7
tmp(325) := SUB & REG_7 & "0000000111"; --  Decrementa o valor das dezenas dos minutos do timer
tmp(326) := STA & REG_7 & "0000011000"; --  Salva o valor das dezenas dos minutos do timer
tmp(327) := LDA & REG_7 & "0000100011"; --  Carrega o valor -1 para R7
tmp(328) := CHECK & REG_7 & "0000011000"; --  Verifica se o valor das dezenas dos minutos do timer é igual a -1
tmp(329) := JNE & REG_0 & "1001100001"; -- JNE
tmp(330) := LDI & REG_3 & "0000000101"; --  Seta o valor 5 para R3
tmp(331) := STA & REG_3 & "0000011000"; --  Salva o valor 5 nas dezenas dos minutos do timer
tmp(332) := LDA & REG_7 & "0000011001"; --  Carrega o valor das unidades das horas do timer para R7
tmp(333) := SUB & REG_7 & "0000000111"; --  Decrementa o valor das unidades das horas do timer
tmp(334) := STA & REG_7 & "0000011001"; --  Salva o valor das unidades das horas do timer
tmp(335) := LDA & REG_7 & "0000100011"; --  Carrega o valor -1 para R7
tmp(336) := CHECK & REG_7 & "0000011001"; --  Verifica se o valor das unidades das horas do timer é igual a -1
tmp(337) := JNE & REG_0 & "1001100001"; -- JNE
tmp(338) := LDI & REG_3 & "0000001001"; --  Seta o valor 9 para R3
tmp(339) := STA & REG_3 & "0000011001"; --  Salva o valor 9 nas unidades das horas do timer
tmp(340) := LDA & REG_7 & "0000011010"; --  Carrega o valor das dezenas das horas do timer para R7
tmp(341) := SUB & REG_7 & "0000000111"; --  Decrementa o valor das dezenas das horas do timer
tmp(342) := STA & REG_7 & "0000011010"; --  Salva o valor das dezenas das horas do timer
tmp(343) := LDA & REG_7 & "0000100011"; --  Carrega o valor -1 para R7
tmp(344) := CHECK & REG_7 & "0000011010"; --  Verifica se o valor das dezenas das horas do timer é igual a -1
tmp(345) := JNE & REG_0 & "1001100001"; -- JNE
tmp(346) := STA & REG_1 & "0000100100"; --  Ativa a flag de timer finalizado
tmp(347) := STA & REG_0 & "0000011011"; --  Desativa a flag de timer
tmp(348) := STA & REG_0 & "0000010101"; --  0 -> Novo valor das unidades dos segundos
tmp(349) := STA & REG_0 & "0000010110"; --  0 -> Novo valor das dezenas dos segundos
tmp(350) := STA & REG_0 & "0000010111"; --  0 -> Novo valor das unidades dos minutos
tmp(351) := STA & REG_0 & "0000011000"; --  0 -> Novo valor das dezenas dos minutos
tmp(352) := STA & REG_0 & "0000011001"; --  0 -> Novo valor das unidades das horas
tmp(353) := STA & REG_0 & "0000011010"; --  0 -> Novo valor das dezenas das horas
tmp(354) := STA & REG_0 & "0000011100"; --  Desativa a flag de ajuste das unidades dos segundos do timer
tmp(355) := STA & REG_0 & "0000011101"; --  Desativa a flag de ajuste das dezenas dos segundos do timer
tmp(356) := STA & REG_0 & "0000011110"; --  Desativa a flag de ajuste das unidades dos minutos do timer
tmp(357) := STA & REG_0 & "0000011111"; --  Desativa a flag de ajuste das dezenas dos minutos do timer
tmp(358) := STA & REG_0 & "0000100000"; --  Desativa a flag de ajuste das unidades das horas do timer
tmp(359) := STA & REG_0 & "0000100001"; --  Desativa a flag de ajuste das dezenas (>= 2) das horas do timer
tmp(360) := STA & REG_0 & "0000100010"; --  Desativa a flag de ajuste das dezenas (< 2) das horas do timer
tmp(361) := STA & REG_0 & "0100000000"; --  Apaga os LEDR0 até LEDR7
tmp(362) := STA & REG_0 & "0100000001"; --  Apaga o LEDR8
tmp(363) := RET & REG_0 & "0000000000"; -- RET
tmp(364) := LDA & REG_7 & "0101100011"; --  Carrega o valor do botão KEY3
tmp(365) := ANDI & REG_7 & "0000000111"; --  Aplica máscara AND para isolar o bit 0
tmp(366) := CHECK & REG_7 & "0000000111"; --  Se KEY1 estiver pressionada, passa a setar o limite de incremento
tmp(367) := STA & REG_0 & "0111111100"; -- STA
tmp(368) := JNE & REG_0 & "1001100001"; -- JNE
tmp(369) := LDA & REG_7 & "0000000101"; --  Carrega o valor das dezenas das horas para R7
tmp(370) := CHECK & REG_7 & "0000001010"; --  Verifica se o valor das dezenas das horas é menor que 2
tmp(371) := JLT & REG_0 & "0101111101"; -- JLT
tmp(372) := LDA & REG_7 & "0000000100"; --  Carrega o valor das unidades das horas para R7
tmp(373) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das unidades das horas
tmp(374) := STA & REG_7 & "0000000100"; --  Salva o valor das unidades das horas
tmp(375) := LDA & REG_7 & "0000000100"; --  Carrega o valor das unidades das horas para R7
tmp(376) := CHECK & REG_7 & "0000001011"; --  Verifica se o valor das unidades das horas é menor que 4
tmp(377) := JLT & REG_0 & "1001100001"; -- JLT
tmp(378) := STA & REG_0 & "0000000100"; --  0 -> Valor das unidades das horas
tmp(379) := STA & REG_0 & "0000000101"; --  0 -> Valor das dezenas das horas
tmp(380) := RET & REG_0 & "0000000000"; -- RET
tmp(381) := LDA & REG_7 & "0000000100"; --  Carrega o valor das unidades das horas para R7
tmp(382) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das unidades das horas
tmp(383) := STA & REG_7 & "0000000100"; --  Salva o valor das unidades das horas
tmp(384) := LDA & REG_7 & "0000000100"; --  Carrega o valor das unidades das horas para R7
tmp(385) := CHECK & REG_7 & "0000001000"; --  Verifica se o valor das unidades das horas é menor que 10
tmp(386) := JLT & REG_0 & "1001100001"; -- JLT
tmp(387) := STA & REG_0 & "0000000100"; --  0 -> Valor das unidades das horas
tmp(388) := LDA & REG_7 & "0000000101"; --  Carrega o valor das dezenas das horas para R7
tmp(389) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das dezenas das horas
tmp(390) := STA & REG_7 & "0000000101"; --  Salva o valor das dezenas das horas
tmp(391) := RET & REG_0 & "0000000000"; -- RET
tmp(392) := LDA & REG_7 & "0101100010"; --  Carrega o valor do botão KEY2
tmp(393) := ANDI & REG_7 & "0000000111"; --  Aplica máscara AND para isolar o bit 0
tmp(394) := CHECK & REG_7 & "0000000111"; --  Se KEY2 estiver pressionada, passa a setar o limite de incremento
tmp(395) := STA & REG_0 & "0111111101"; -- STA
tmp(396) := JNE & REG_0 & "1001100001"; -- JNE
tmp(397) := LDA & REG_7 & "0000000010"; --  Carrega o valor das unidades dos minutos para R7
tmp(398) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das unidades dos minutos
tmp(399) := STA & REG_7 & "0000000010"; --  Salva o valor das unidades dos minutos
tmp(400) := LDA & REG_7 & "0000000010"; --  Carrega o valor das unidades dos minutos para R7
tmp(401) := CHECK & REG_7 & "0000001000"; --  Verifica se o valor das unidades dos minutos é menor que 10
tmp(402) := JLT & REG_0 & "1001100001"; -- JLT
tmp(403) := STA & REG_0 & "0000000010"; --  0 -> Valor das unidades dos minutos
tmp(404) := LDA & REG_7 & "0000000011"; --  Carrega o valor das dezenas dos minutos para R7
tmp(405) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das dezenas dos minutos
tmp(406) := STA & REG_7 & "0000000011"; --  Salva o valor das dezenas dos minutos
tmp(407) := LDA & REG_7 & "0000000011"; --  Carrega o valor das dezenas dos minutos para R7
tmp(408) := CHECK & REG_7 & "0000001001"; --  Verifica se o valor das dezenas dos minutos é menor que 6
tmp(409) := JLT & REG_0 & "1001100001"; -- JLT
tmp(410) := STA & REG_0 & "0000000011"; --  0 -> Valor das dezenas dos minutos
tmp(411) := RET & REG_0 & "0000000000"; -- RET
tmp(412) := LDA & REG_7 & "0101100001"; --  Carrega o valor do botão KEY1
tmp(413) := ANDI & REG_7 & "0000000111"; --  Aplica máscara AND para isolar o bit 0
tmp(414) := CHECK & REG_7 & "0000000111"; --  Se KEY1 estiver pressionada, passa a setar o limite de incremento
tmp(415) := STA & REG_0 & "0111111110"; -- STA
tmp(416) := JNE & REG_0 & "1001100001"; -- JNE
tmp(417) := LDA & REG_7 & "0000000000"; --  Carrega o valor das unidades dos segundos para R7
tmp(418) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das unidades dos segundos
tmp(419) := STA & REG_7 & "0000000000"; --  Salva o valor das unidades dos segundos
tmp(420) := LDA & REG_7 & "0000000000"; --  Carrega o valor das unidades dos segundos para R7
tmp(421) := CHECK & REG_7 & "0000001000"; --  Verifica se o valor das unidades dos segundos é menor que 10
tmp(422) := JLT & REG_0 & "1001100001"; -- JLT
tmp(423) := STA & REG_0 & "0000000000"; --  0 -> Valor das unidades dos segundos
tmp(424) := LDA & REG_7 & "0000000001"; --  Carrega o valor das dezenas dos segundos para R7
tmp(425) := SOMA & REG_7 & "0000000111"; --  Incrementa o valor das dezenas dos segundos
tmp(426) := STA & REG_7 & "0000000001"; --  Salva o valor das dezenas dos segundos
tmp(427) := LDA & REG_7 & "0000000001"; --  Carrega o valor das dezenas dos segundos para R7
tmp(428) := CHECK & REG_7 & "0000001001"; --  Verifica se o valor das dezenas dos segundos é menor que 6
tmp(429) := JLT & REG_0 & "1001100001"; -- JLT
tmp(430) := STA & REG_0 & "0000000001"; --  0 -> Valor das dezenas dos segundos
tmp(431) := RET & REG_0 & "0000000000"; -- RET
tmp(432) := LDA & REG_7 & "0101000000"; --  Carrega o R7 com a leitura das chaves SW0 até SW7
tmp(433) := ANDI & REG_7 & "0000001100"; --  Aplica máscara AND para isolar o bit 7
tmp(434) := CHECK & REG_7 & "0000001100"; --  Verifica se a chave SW7 está pressionada
tmp(435) := JNE & REG_0 & "1001100001"; -- JNE
tmp(436) := LDA & REG_7 & "0101100000"; --  Carrega o valor do botão KEY0
tmp(437) := ANDI & REG_7 & "0000000111"; --  Aplica máscara AND para isolar o bit 0
tmp(438) := CHECK & REG_7 & "0000000111"; --  Se KEY0 estiver pressionada, passa a setar o limite de incremento
tmp(439) := STA & REG_0 & "0111111111"; -- STA
tmp(440) := JNE & REG_0 & "1001100001"; -- JNE
tmp(441) := LDA & REG_7 & "0000001110"; --  Carrega o valor da flag de alarme para R7
tmp(442) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de alarme está setada
tmp(443) := JEQ & REG_0 & "1001100001"; -- JEQ
tmp(444) := JSR & REG_0 & "1001010101"; -- JSR
tmp(445) := STA & REG_1 & "0100000010"; --  Acende o LEDR9 para indicar que é o alarme que está sendo setado
tmp(446) := LDA & REG_7 & "0000101011"; --  Carrega o valor da flag de ajuste das dezenas (< 2) das horas para R7
tmp(447) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das dezenas das horas está setada
tmp(448) := JEQ & REG_0 & "0111010000"; -- JEQ
tmp(449) := LDA & REG_7 & "0000101010"; --  Carrega o valor da flag de ajuste das dezenas (>= 2) das horas para R7
tmp(450) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das dezenas das horas está setada
tmp(451) := JEQ & REG_0 & "0111011111"; -- JEQ
tmp(452) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(453) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(454) := STA & REG_7 & "0000010100"; --  Salva o valor de SW0 até SW7 em @20
tmp(455) := LDA & REG_7 & "0000010100"; --  Carrega o valor de SW0 até SW7 para R7
tmp(456) := CHECK & REG_7 & "0000001010"; --  Compara o valor de SW0 até SW7 com 2
tmp(457) := JLT & REG_0 & "0111001100"; -- JLT
tmp(458) := JEQ & REG_0 & "0111011010"; -- JEQ
tmp(459) := JMP & REG_0 & "1001100001"; -- JMP
tmp(460) := LDI & REG_3 & "0000100000"; --  Seta o valor 32 para R3
tmp(461) := STA & REG_3 & "0100000000"; --  Acende o LEDR5 para indicar que o valor das dezenas das horas do alarme foi setado
tmp(462) := STA & REG_1 & "0000101011"; --  Ativa a flag de ajuste das dezenas das horas
tmp(463) := RET & REG_0 & "0000000000"; -- RET
tmp(464) := LDA & REG_7 & "0000101001"; --  Carrega o valor da flag de ajuste das unidades das horas para R7
tmp(465) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das unidades das horas está setada
tmp(466) := JEQ & REG_0 & "0111101110"; -- JEQ
tmp(467) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(468) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(469) := STA & REG_7 & "0000010011"; --  Salva o valor de SW0 até SW7 em @19
tmp(470) := LDA & REG_7 & "0000010011"; --  Carrega o valor de SW0 até SW7 para R7
tmp(471) := CHECK & REG_7 & "0000001000"; --  Compara o valor de SW0 até SW7 com 10
tmp(472) := JLT & REG_0 & "0111101001"; -- JLT
tmp(473) := JMP & REG_0 & "1001100001"; -- JMP
tmp(474) := LDI & REG_3 & "0000100000"; --  Seta o valor 32 para R3
tmp(475) := STA & REG_3 & "0100000000"; --  Acende o LEDR5 para indicar que o valor das dezenas das horas do alarme foi setado
tmp(476) := STA & REG_1 & "0000101010"; --  Ativa a flag de ajuste das dezenas das horas
tmp(477) := STA & REG_1 & "0100000010"; --  Acende o LEDR9 para indicar que é o alarme que está sendo setado, e não o timer
tmp(478) := RET & REG_0 & "0000000000"; -- RET
tmp(479) := LDA & REG_7 & "0000101001"; --  Carrega o valor da flag de ajuste das unidades das horas para R7
tmp(480) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das unidades das horas está setada
tmp(481) := JEQ & REG_0 & "0111101110"; -- JEQ
tmp(482) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(483) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(484) := STA & REG_7 & "0000010011"; --  Salva o valor de SW0 até SW7 em @19
tmp(485) := LDA & REG_7 & "0000010011"; --  Carrega o valor de SW0 até SW7 para R7
tmp(486) := CHECK & REG_7 & "0000001011"; --  Compara o valor de SW0 até SW7 com 4
tmp(487) := JLT & REG_0 & "0111101001"; -- JLT
tmp(488) := JMP & REG_0 & "1001100001"; -- JMP
tmp(489) := LDI & REG_3 & "0000110000"; --  Seta o valor 48 para R3
tmp(490) := STA & REG_3 & "0100000000"; --  Acende o LEDR5 e LEDR4 para indicar que os valores das dezenas e unidade de horas do alarme foram setados
tmp(491) := STA & REG_1 & "0000101001"; --  Ativa a flag de ajuste das unidades das horas
tmp(492) := STA & REG_1 & "0100000010"; --  Acende o LEDR9 para indicar que é o alarme que está sendo setado, e não o timer
tmp(493) := RET & REG_0 & "0000000000"; -- RET
tmp(494) := LDA & REG_7 & "0000101000"; --  Carrega o valor da flag de ajuste das dezenas dos minutos para R7
tmp(495) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das dezenas dos minutos está setada
tmp(496) := JEQ & REG_0 & "0111111101"; -- JEQ
tmp(497) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(498) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(499) := STA & REG_7 & "0000010010"; --  Salva o valor de SW0 até SW7 em @18
tmp(500) := LDA & REG_7 & "0000010010"; --  Carrega o valor de SW0 até SW7 para R7
tmp(501) := CHECK & REG_7 & "0000001001"; --  Compara o valor de SW0 até SW7 com 6
tmp(502) := JLT & REG_0 & "0111111000"; -- JLT
tmp(503) := JMP & REG_0 & "1001100001"; -- JMP
tmp(504) := LDI & REG_3 & "0000111000"; --  Seta o valor 56 para R3
tmp(505) := STA & REG_3 & "0100000000"; --  Acende o LEDR5, LEDR4 e LEDR3 para indicar que os valores das dezenas, unidade de horas e dezenas de minutos do alarme foram setados
tmp(506) := STA & REG_1 & "0000101000"; --  Ativa a flag de ajuste das dezenas dos minutos
tmp(507) := STA & REG_1 & "0100000010"; --  Acende o LEDR9 para indicar que é o alarme que está sendo setado, e não o timer
tmp(508) := RET & REG_0 & "0000000000"; -- RET
tmp(509) := LDA & REG_7 & "0000100111"; --  Carrega o valor da flag de ajuste das unidades dos minutos para R7
tmp(510) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das unidades dos minutos está setada
tmp(511) := JEQ & REG_0 & "1000001100"; -- JEQ
tmp(512) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(513) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(514) := STA & REG_7 & "0000010001"; --  Salva o valor de SW0 até SW7 em @17
tmp(515) := LDA & REG_7 & "0000010001"; --  Carrega o valor de SW0 até SW7 para R7
tmp(516) := CHECK & REG_7 & "0000001000"; --  Compara o valor de SW0 até SW7 com 10
tmp(517) := JLT & REG_0 & "1000000111"; -- JLT
tmp(518) := JMP & REG_0 & "1001100001"; -- JMP
tmp(519) := LDI & REG_3 & "0000111100"; --  Seta o valor 60 para R3
tmp(520) := STA & REG_3 & "0100000000"; --  Acende os LEDR5, LEDR4, LEDR3 e LEDR2 para indicar que os valores das dezenas, unidade de horas e dezenas de minutos do alarme foram setados
tmp(521) := STA & REG_1 & "0000100111"; --  Ativa a flag de ajuste das unidades dos minutos
tmp(522) := STA & REG_1 & "0100000010"; --  Acende o LEDR9 para indicar que é o alarme que está sendo setado, e não o timer
tmp(523) := RET & REG_0 & "0000000000"; -- RET
tmp(524) := LDA & REG_7 & "0000100110"; --  Carrega o valor da flag de ajuste das dezenas dos segundos para R7
tmp(525) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das dezenas dos segundos está setada
tmp(526) := JEQ & REG_0 & "1000011011"; -- JEQ
tmp(527) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(528) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(529) := STA & REG_7 & "0000010000"; --  Salva o valor de SW0 até SW7 em @16
tmp(530) := LDA & REG_7 & "0000010000"; --  Carrega o valor de SW0 até SW7 para R7
tmp(531) := CHECK & REG_7 & "0000001001"; --  Compara o valor de SW0 até SW7 com 6
tmp(532) := JLT & REG_0 & "1000010110"; -- JLT
tmp(533) := JMP & REG_0 & "1001100001"; -- JMP
tmp(534) := LDI & REG_3 & "0000111110"; --  Seta o valor 62 para R3
tmp(535) := STA & REG_3 & "0100000000"; --  Acende o LEDR5, LEDR4, LEDR3, LEDR2 e LEDR1 para indicar que os valores das dezenas, unidade de horas, dezenas e unidade dos minutos do alarme foram setados
tmp(536) := STA & REG_1 & "0000100110"; --  Ativa a flag de ajuste das dezenas dos segundos
tmp(537) := STA & REG_1 & "0100000010"; --  Acende o LEDR9 para indicar que é o alarme que está sendo setado, e não o timer
tmp(538) := RET & REG_0 & "0000000000"; -- RET
tmp(539) := LDA & REG_7 & "0000100101"; --  Carrega o valor da flag de ajuste das unidades dos segundos para R7
tmp(540) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de ajuste das unidades dos segundos está setada
tmp(541) := JEQ & REG_0 & "1000100101"; -- JEQ
tmp(542) := LDA & REG_7 & "0101000000"; --  Carrega o r7 com a leitura das chaves SW0 até SW7
tmp(543) := ANDI & REG_7 & "0000101101"; --  Aplica máscara AND para não haver leitura do SW7 ~ SW4
tmp(544) := STA & REG_7 & "0000001111"; --  Salva o valor de SW0 até SW7 em @15
tmp(545) := LDA & REG_7 & "0000001111"; --  Carrega o valor de SW0 até SW7 para R7
tmp(546) := CHECK & REG_7 & "0000001000"; --  Compara o valor de SW0 até SW7 com 10
tmp(547) := JLT & REG_0 & "1000100101"; -- JLT
tmp(548) := JMP & REG_0 & "1001100001"; -- JMP
tmp(549) := LDI & REG_3 & "0000111111"; --  Seta o valor 63 para R3
tmp(550) := STA & REG_3 & "0100000000"; --  Acende o LEDR5, LEDR4, LEDR3, LEDR2, LEDR1 e LEDR0 para indicar que os valores das dezenas, unidade de horas, dezenas e unidade de minutos e dezenas e unidade dos segundos do alarme foram setados
tmp(551) := STA & REG_1 & "0000001110"; --  Ativa a flag de alarme setado
tmp(552) := RET & REG_0 & "0000000000"; -- RET
tmp(553) := LDA & REG_7 & "0000101100"; --  Carrega o valor da flag de alarme atingido para R7
tmp(554) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de alarme atingido está setada
tmp(555) := JEQ & REG_0 & "1001000011"; -- JEQ
tmp(556) := LDA & REG_7 & "0000001110"; --  Carrega o valor da flag de alarme setado para R7
tmp(557) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de alarme setado está setada
tmp(558) := JNE & REG_0 & "1001100001"; -- JNE
tmp(559) := LDA & REG_7 & "0000000101"; --  Carrega o valor das dezenas das horas do alarme para R7
tmp(560) := CHECK & REG_7 & "0000010100"; --  Verifica se o valor das dezenas das horas do alarme é igual ao valor das dezenas das horas do timer
tmp(561) := JNE & REG_0 & "1001100001"; -- JNE
tmp(562) := LDA & REG_7 & "0000000100"; --  Carrega o valor das unidades das horas do alarme para R7
tmp(563) := CHECK & REG_7 & "0000010011"; --  Verifica se o valor das unidades das horas do alarme é igual ao valor das unidades das horas do timer
tmp(564) := JNE & REG_0 & "1001100001"; -- JNE
tmp(565) := LDA & REG_7 & "0000000011"; --  Carrega o valor das dezenas dos minutos do alarme para R7
tmp(566) := CHECK & REG_7 & "0000010010"; --  Verifica se o valor das dezenas dos minutos do alarme é igual ao valor das dezenas dos minutos do timer
tmp(567) := JNE & REG_0 & "1001100001"; -- JNE
tmp(568) := LDA & REG_7 & "0000000010"; --  Carrega o valor das unidades dos minutos do alarme para R7
tmp(569) := CHECK & REG_7 & "0000010001"; --  Verifica se o valor das unidades dos minutos do alarme é igual ao valor das unidades dos minutos do timer
tmp(570) := JNE & REG_0 & "1001100001"; -- JNE
tmp(571) := LDA & REG_7 & "0000000001"; --  Carrega o valor das dezenas dos segundos do alarme para R7
tmp(572) := CHECK & REG_7 & "0000010000"; --  Verifica se o valor das dezenas dos segundos do alarme é igual ao valor das dezenas dos segundos do timer
tmp(573) := JNE & REG_0 & "1001100001"; -- JNE
tmp(574) := LDA & REG_7 & "0000000000"; --  Carrega o valor das unidades dos segundos do alarme para R7
tmp(575) := CHECK & REG_7 & "0000001111"; --  Verifica se o valor das unidades dos segundos do alarme é igual ao valor das unidades dos segundos do timer
tmp(576) := JNE & REG_0 & "1001100001"; -- JNE
tmp(577) := STA & REG_1 & "0000101100"; --  Ativa a flag de alarme atingido
tmp(578) := RET & REG_0 & "0000000000"; -- RET
tmp(579) := STA & REG_0 & "0100000010"; --  Apaga o LEDR9 para indicar que o alarme foi atingido
tmp(580) := STA & REG_0 & "0100000000"; --  Apaga os LEDs de ajuste e valor do alarme
tmp(581) := STA & REG_0 & "0000001110"; --  0 -> Flag de alarme setado
tmp(582) := STA & REG_0 & "0000001111"; --  0 -> Valor das unidades dos segundos do alarme
tmp(583) := STA & REG_0 & "0000010000"; --  0 -> Valor das dezenas dos segundos do alarme
tmp(584) := STA & REG_0 & "0000010001"; --  0 -> Valor das unidades dos minutos do alarme
tmp(585) := STA & REG_0 & "0000010010"; --  0 -> Valor das dezenas dos minutos do alarme
tmp(586) := STA & REG_0 & "0000010011"; --  0 -> Valor das unidades das horas do alarme
tmp(587) := STA & REG_0 & "0000010100"; --  0 -> Valor das dezenas das horas do alarme
tmp(588) := STA & REG_0 & "0000100101"; --  0 -> Flag de ajuste das unidades dos segundos do alarme
tmp(589) := STA & REG_0 & "0000100110"; --  0 -> Flag de ajuste das dezenas dos segundos
tmp(590) := STA & REG_0 & "0000100111"; --  0 -> Flag de ajuste das unidades dos segundos
tmp(591) := STA & REG_0 & "0000101000"; --  0 -> Flag de ajuste das dezenas dos minutos
tmp(592) := STA & REG_0 & "0000101001"; --  0 -> Flag de ajuste das unidades dos minutos
tmp(593) := STA & REG_0 & "0000101010"; --  0 -> Flag de ajuste das dezenas (>= 2) das horas
tmp(594) := STA & REG_0 & "0000101011"; --  0 -> Flag de ajuste das dezenas (< 2) das horas
tmp(595) := STA & REG_0 & "0000101100"; --  0 -> Flag de chegou no horário do alarme
tmp(596) := RET & REG_0 & "0000000000"; -- RET
tmp(597) := STA & REG_0 & "0100000001"; --  Apaga o LEDR8
tmp(598) := LDA & REG_7 & "0000011011"; --  Carrega o valor da flag de timer setado para R7
tmp(599) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de timer setado está setada
tmp(600) := JNE & REG_0 & "1001100001"; -- JNE
tmp(601) := STA & REG_1 & "0100000001"; --  Acende o LEDR8
tmp(602) := RET & REG_0 & "0000000000"; -- RET
tmp(603) := STA & REG_0 & "0100000010"; --  Apaga o LEDR9
tmp(604) := LDA & REG_7 & "0000001110"; --  Carrega o valor da flag de alarme setado para R7
tmp(605) := CHECK & REG_7 & "0000000111"; --  Verifica se a flag de alarme setado está setada
tmp(606) := JNE & REG_0 & "1001100001"; -- JNE
tmp(607) := STA & REG_1 & "0100000010"; --  Acende o LEDR9
tmp(608) := RET & REG_0 & "0000000000"; -- RET
tmp(609) := RET & REG_0 & "0000000000"; -- RET

		  return tmp;
    end initMemory;


  -- Sinal que armazena os dados da função initMemory.
  signal memROM : blocoMemoria := initMemory;

begin
  -- Saída de dados baseada no endereço de entrada.
  Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;